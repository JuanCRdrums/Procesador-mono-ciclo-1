
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity RF is
    port (
          RD : in std_logic_vector(4 downto 0);
          DWR   : in std_logic_vector(31 downto 0);
			 RS1   : in std_logic_vector(4 downto 0);
			 RS2   : in std_logic_vector(4 downto 0);
          CRS1   : out std_logic_vector(31 downto 0);
			 CRS2   : out std_logic_vector(31 downto 0);
			 rst: in std_logic
			 );
end RF;

architecture syn of RF is
    type ram_type is array (0 to 31) of std_logic_vector (31 downto 0);
    signal RAM: ram_type;
begin

    process (RD,DWR,RS1,RS2,rst)
    begin
			RAM(0) <= "00000000000000000000000000000000";
			CRS1 <= RAM(conv_integer(RS1));
			CRS2 <= RAM(conv_integer(RS2));
			if(RD /= "00000") then
				RAM(conv_integer(RD)) <= DWR;
			end if;
        if rst = '1' then
				RAM(0) <= "00000000000000000000000000000000";
				RAM(1) <= "00000000000000000000000000000000";
				RAM(2) <= "00000000000000000000000000000000";
				RAM(3) <= "00000000000000000000000000000000";
				RAM(4) <= "00000000000000000000000000000000";
				RAM(5) <= "00000000000000000000000000000000";
				RAM(6) <= "00000000000000000000000000000000";
				RAM(7) <= "00000000000000000000000000000000";
				RAM(8) <= "00000000000000000000000000000000";
				RAM(9) <= "00000000000000000000000000000000";
				RAM(10) <= "00000000000000000000000000000000";
				RAM(11) <= "00000000000000000000000000000000";
				RAM(12) <= "00000000000000000000000000000000";
				RAM(13) <= "00000000000000000000000000000000";
				RAM(14) <= "00000000000000000000000000000000";
				RAM(15) <= "00000000000000000000000000000000";
				RAM(16) <= "00000000000000000000000000000000";
				RAM(17) <= "00000000000000000000000000000000";
				RAM(18) <= "00000000000000000000000000000000";
				RAM(19) <= "00000000000000000000000000000000";
				RAM(20) <= "00000000000000000000000000000000";
				RAM(21) <= "00000000000000000000000000000000";
				RAM(22) <= "00000000000000000000000000000000";
				RAM(23) <= "00000000000000000000000000000000";
				RAM(24) <= "00000000000000000000000000000000";
				RAM(25) <= "00000000000000000000000000000000";
				RAM(26) <= "00000000000000000000000000000000";
				RAM(27) <= "00000000000000000000000000000000";
				RAM(28) <= "00000000000000000000000000000000";
				RAM(29) <= "00000000000000000000000000000000";
				RAM(30) <= "00000000000000000000000000000000";
				RAM(31) <= "00000000000000000000000000000000";				
        end if;
    end process;

end syn;